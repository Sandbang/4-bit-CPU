`timescale 1ns / 1ps

module main_tb();


endmodule
